library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

ENTITY main IS
	
PORT(a,b,c:IN std_logic;
d: OUT std_logic);

END main;

ARCHITECTURE myMain OF main IS
BEGIN

END myMain;