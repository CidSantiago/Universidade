LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY mux16x1 IS 

PORT (
